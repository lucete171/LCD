//testbench of computation_1

//timescale `timescale 1ns/1ns
module tb_sm;
  PE_module PE_1(.A(), .B(), 
  
  
endmodule